// modulo decodificacion de la tecla presionada del teclado
module decoder_keyb(
    input wire key_coord[0:7],
    input wire button_pressed,
    output wire key[0:1],
    input wire clk
);

assign 

always @(posedge clk) begin
    if (button_pressed) 
end
endmodule