// main
module top (
    ports sape
);
    
endmodule